RAIZQUADRADA_inst : RAIZQUADRADA PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		result	 => result_sig
	);
