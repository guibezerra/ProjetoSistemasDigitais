Constante2_inst : Constante2 PORT MAP (
		result	 => result_sig
	);
