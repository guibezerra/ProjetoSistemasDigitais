EXP1_inst : EXP1 PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		result	 => result_sig
	);
