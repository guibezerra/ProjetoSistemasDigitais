Constante_0_inst : Constante_0 PORT MAP (
		result	 => result_sig
	);
