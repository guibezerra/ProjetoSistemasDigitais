-- megafunction wizard: %ALTFP_CONVERT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTFP_CONVERT 

-- ============================================================
-- File Name: ConvIntToFloat.vhd
-- Megafunction Name(s):
-- 			ALTFP_CONVERT
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 17.1.0 Build 590 10/25/2017 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2017  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details.


--altfp_convert CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" OPERATION="INT2FLOAT" ROUNDING="TO_NEAREST" WIDTH_DATA=10 WIDTH_EXP_INPUT=8 WIDTH_EXP_OUTPUT=8 WIDTH_INT=10 WIDTH_MAN_INPUT=23 WIDTH_MAN_OUTPUT=23 WIDTH_RESULT=32 clock dataa result
--VERSION_BEGIN 17.1 cbx_altbarrel_shift 2017:10:25:18:06:52:SJ cbx_altera_syncram_nd_impl 2017:10:25:18:06:52:SJ cbx_altfp_convert 2017:10:25:18:06:52:SJ cbx_altpriority_encoder 2017:10:25:18:06:52:SJ cbx_altsyncram 2017:10:25:18:06:53:SJ cbx_cycloneii 2017:10:25:18:06:53:SJ cbx_lpm_abs 2017:10:25:18:06:53:SJ cbx_lpm_add_sub 2017:10:25:18:06:53:SJ cbx_lpm_compare 2017:10:25:18:06:53:SJ cbx_lpm_decode 2017:10:25:18:06:53:SJ cbx_lpm_divide 2017:10:25:18:06:53:SJ cbx_lpm_mux 2017:10:25:18:06:53:SJ cbx_mgl 2017:10:25:18:08:29:SJ cbx_nadder 2017:10:25:18:06:53:SJ cbx_stratix 2017:10:25:18:06:53:SJ cbx_stratixii 2017:10:25:18:06:53:SJ cbx_stratixiii 2017:10:25:18:06:53:SJ cbx_stratixv 2017:10:25:18:06:53:SJ cbx_util_mgl 2017:10:25:18:06:53:SJ  VERSION_END


--altbarrel_shift CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" PIPELINE=2 SHIFTDIR="LEFT" SHIFTTYPE="LOGICAL" WIDTH=10 WIDTHDIST=4 aclr clk_en clock data distance result
--VERSION_BEGIN 17.1 cbx_altbarrel_shift 2017:10:25:18:06:52:SJ cbx_mgl 2017:10:25:18:08:29:SJ  VERSION_END

--synthesis_resources = reg 24 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  ConvIntToFloat_altbarrel_shift_aof IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clk_en	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (9 DOWNTO 0);
		 distance	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (9 DOWNTO 0)
	 ); 
 END ConvIntToFloat_altbarrel_shift_aof;

 ARCHITECTURE RTL OF ConvIntToFloat_altbarrel_shift_aof IS

	 SIGNAL	 dir_pipe	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper1d	:	STD_LOGIC_VECTOR(9 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper2d	:	STD_LOGIC_VECTOR(9 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec2r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec3r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range46w58w59w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range46w54w55w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range67w79w80w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range67w75w76w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range90w101w102w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range90w97w98w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range109w120w121w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range109w116w117w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range46w50w51w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range67w71w72w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range90w93w94w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range109w112w113w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range46w58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range46w54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range67w79w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range67w75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range90w101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range90w97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range109w120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range109w116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range43w57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range65w78w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range88w100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range107w119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range46w50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range67w71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range90w93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range109w112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range46w58w59w60w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range67w79w80w81w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range90w101w102w103w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range109w120w121w122w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_lg_w_sel_w_range46w58w59w60w61w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_lg_w_sel_w_range67w79w80w81w82w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w104w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w123w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  dir_w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  direction_w :	STD_LOGIC;
	 SIGNAL  pad_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  sbit_w :	STD_LOGIC_VECTOR (49 DOWNTO 0);
	 SIGNAL  sel_w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  smux_w :	STD_LOGIC_VECTOR (39 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w115w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w118w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_w_pad_w_range48w_w_w_sbit_w_range41w_range52w53w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_w_pad_w_range69w_w_w_sbit_w_range64w_range73w74w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_w_pad_w_range91w_w_w_sbit_w_range84w_range95w96w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_w_w_sbit_w_range41w_range49w_w_pad_w_range48w56w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_w_w_sbit_w_range64w_range70w_w_pad_w_range69w77w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_w_w_sbit_w_range84w_range92w_w_pad_w_range91w99w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range43w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range88w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range64w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range84w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range106w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range41w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range46w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_smux_w_range83w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_smux_w_range124w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
 BEGIN

	loop0 : FOR i IN 0 TO 9 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range46w58w59w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range46w58w(0) AND wire_altbarrel_shift5_w_w_w_sbit_w_range41w_range49w_w_pad_w_range48w56w(i);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 9 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range46w54w55w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range46w54w(0) AND wire_altbarrel_shift5_w_w_pad_w_range48w_w_w_sbit_w_range41w_range52w53w(i);
	END GENERATE loop1;
	loop2 : FOR i IN 0 TO 9 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range67w79w80w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range67w79w(0) AND wire_altbarrel_shift5_w_w_w_sbit_w_range64w_range70w_w_pad_w_range69w77w(i);
	END GENERATE loop2;
	loop3 : FOR i IN 0 TO 9 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range67w75w76w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range67w75w(0) AND wire_altbarrel_shift5_w_w_pad_w_range69w_w_w_sbit_w_range64w_range73w74w(i);
	END GENERATE loop3;
	loop4 : FOR i IN 0 TO 9 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range90w101w102w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range90w101w(0) AND wire_altbarrel_shift5_w_w_w_sbit_w_range84w_range92w_w_pad_w_range91w99w(i);
	END GENERATE loop4;
	loop5 : FOR i IN 0 TO 9 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range90w97w98w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range90w97w(0) AND wire_altbarrel_shift5_w_w_pad_w_range91w_w_w_sbit_w_range84w_range95w96w(i);
	END GENERATE loop5;
	loop6 : FOR i IN 0 TO 9 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range109w120w121w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range109w120w(0) AND wire_altbarrel_shift5_w118w(i);
	END GENERATE loop6;
	loop7 : FOR i IN 0 TO 9 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range109w116w117w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range109w116w(0) AND wire_altbarrel_shift5_w115w(i);
	END GENERATE loop7;
	loop8 : FOR i IN 0 TO 9 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range46w50w51w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range46w50w(0) AND wire_altbarrel_shift5_w_sbit_w_range41w(i);
	END GENERATE loop8;
	loop9 : FOR i IN 0 TO 9 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range67w71w72w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range67w71w(0) AND wire_altbarrel_shift5_w_sbit_w_range64w(i);
	END GENERATE loop9;
	loop10 : FOR i IN 0 TO 9 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range90w93w94w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range90w93w(0) AND wire_altbarrel_shift5_w_sbit_w_range84w(i);
	END GENERATE loop10;
	loop11 : FOR i IN 0 TO 9 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range109w112w113w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range109w112w(0) AND wire_altbarrel_shift5_w_sbit_w_range106w(i);
	END GENERATE loop11;
	wire_altbarrel_shift5_w_lg_w_sel_w_range46w58w(0) <= wire_altbarrel_shift5_w_sel_w_range46w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range43w57w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range46w54w(0) <= wire_altbarrel_shift5_w_sel_w_range46w(0) AND wire_altbarrel_shift5_w_dir_w_range43w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range67w79w(0) <= wire_altbarrel_shift5_w_sel_w_range67w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range65w78w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range67w75w(0) <= wire_altbarrel_shift5_w_sel_w_range67w(0) AND wire_altbarrel_shift5_w_dir_w_range65w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range90w101w(0) <= wire_altbarrel_shift5_w_sel_w_range90w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range88w100w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range90w97w(0) <= wire_altbarrel_shift5_w_sel_w_range90w(0) AND wire_altbarrel_shift5_w_dir_w_range88w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range109w120w(0) <= wire_altbarrel_shift5_w_sel_w_range109w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range107w119w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range109w116w(0) <= wire_altbarrel_shift5_w_sel_w_range109w(0) AND wire_altbarrel_shift5_w_dir_w_range107w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range43w57w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range43w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range65w78w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range65w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range88w100w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range88w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range107w119w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range107w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range46w50w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range46w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range67w71w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range67w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range90w93w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range90w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range109w112w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range109w(0);
	loop12 : FOR i IN 0 TO 9 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range46w58w59w60w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range46w58w59w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range46w54w55w(i);
	END GENERATE loop12;
	loop13 : FOR i IN 0 TO 9 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range67w79w80w81w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range67w79w80w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range67w75w76w(i);
	END GENERATE loop13;
	loop14 : FOR i IN 0 TO 9 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range90w101w102w103w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range90w101w102w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range90w97w98w(i);
	END GENERATE loop14;
	loop15 : FOR i IN 0 TO 9 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range109w120w121w122w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range109w120w121w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range109w116w117w(i);
	END GENERATE loop15;
	loop16 : FOR i IN 0 TO 9 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_lg_w_sel_w_range46w58w59w60w61w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range46w58w59w60w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range46w50w51w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 9 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_lg_w_sel_w_range67w79w80w81w82w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range67w79w80w81w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range67w71w72w(i);
	END GENERATE loop17;
	loop18 : FOR i IN 0 TO 9 GENERATE 
		wire_altbarrel_shift5_w104w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range90w101w102w103w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range90w93w94w(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 9 GENERATE 
		wire_altbarrel_shift5_w123w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range109w120w121w122w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range109w112w113w(i);
	END GENERATE loop19;
	dir_w <= ( dir_pipe(1) & dir_w(2) & dir_pipe(0) & dir_w(0) & direction_w);
	direction_w <= '0';
	pad_w <= (OTHERS => '0');
	result <= sbit_w(49 DOWNTO 40);
	sbit_w <= ( sbit_piper2d & smux_w(29 DOWNTO 20) & sbit_piper1d & smux_w(9 DOWNTO 0) & data);
	sel_w <= ( sel_pipec3r1d & sel_pipec2r1d & distance(1 DOWNTO 0));
	smux_w <= ( wire_altbarrel_shift5_w123w & wire_altbarrel_shift5_w104w & wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_lg_w_sel_w_range67w79w80w81w82w & wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_lg_w_sel_w_range46w58w59w60w61w);
	wire_altbarrel_shift5_w115w <= ( pad_w(7 DOWNTO 0) & sbit_w(39 DOWNTO 38));
	wire_altbarrel_shift5_w118w <= ( sbit_w(31 DOWNTO 30) & pad_w(7 DOWNTO 0));
	wire_altbarrel_shift5_w_w_pad_w_range48w_w_w_sbit_w_range41w_range52w53w <= ( pad_w(0) & sbit_w(9 DOWNTO 1));
	wire_altbarrel_shift5_w_w_pad_w_range69w_w_w_sbit_w_range64w_range73w74w <= ( pad_w(1 DOWNTO 0) & sbit_w(19 DOWNTO 12));
	wire_altbarrel_shift5_w_w_pad_w_range91w_w_w_sbit_w_range84w_range95w96w <= ( pad_w(3 DOWNTO 0) & sbit_w(29 DOWNTO 24));
	wire_altbarrel_shift5_w_w_w_sbit_w_range41w_range49w_w_pad_w_range48w56w <= ( sbit_w(8 DOWNTO 0) & pad_w(0));
	wire_altbarrel_shift5_w_w_w_sbit_w_range64w_range70w_w_pad_w_range69w77w <= ( sbit_w(17 DOWNTO 10) & pad_w(1 DOWNTO 0));
	wire_altbarrel_shift5_w_w_w_sbit_w_range84w_range92w_w_pad_w_range91w99w <= ( sbit_w(25 DOWNTO 20) & pad_w(3 DOWNTO 0));
	wire_altbarrel_shift5_w_dir_w_range43w(0) <= dir_w(0);
	wire_altbarrel_shift5_w_dir_w_range65w(0) <= dir_w(1);
	wire_altbarrel_shift5_w_dir_w_range88w(0) <= dir_w(2);
	wire_altbarrel_shift5_w_dir_w_range107w(0) <= dir_w(3);
	wire_altbarrel_shift5_w_sbit_w_range64w <= sbit_w(19 DOWNTO 10);
	wire_altbarrel_shift5_w_sbit_w_range84w <= sbit_w(29 DOWNTO 20);
	wire_altbarrel_shift5_w_sbit_w_range106w <= sbit_w(39 DOWNTO 30);
	wire_altbarrel_shift5_w_sbit_w_range41w <= sbit_w(9 DOWNTO 0);
	wire_altbarrel_shift5_w_sel_w_range46w(0) <= sel_w(0);
	wire_altbarrel_shift5_w_sel_w_range67w(0) <= sel_w(1);
	wire_altbarrel_shift5_w_sel_w_range90w(0) <= sel_w(2);
	wire_altbarrel_shift5_w_sel_w_range109w(0) <= sel_w(3);
	wire_altbarrel_shift5_w_smux_w_range83w <= smux_w(19 DOWNTO 10);
	wire_altbarrel_shift5_w_smux_w_range124w <= smux_w(39 DOWNTO 30);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dir_pipe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dir_pipe <= ( dir_w(3) & dir_w(1));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper1d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper1d <= wire_altbarrel_shift5_w_smux_w_range83w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper2d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper2d <= wire_altbarrel_shift5_w_smux_w_range124w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec2r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec2r1d <= distance(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec3r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec3r1d <= distance(3);
			END IF;
		END IF;
	END PROCESS;

 END RTL; --ConvIntToFloat_altbarrel_shift_aof


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" WIDTH=16 WIDTHAD=4 data q
--VERSION_BEGIN 17.1 cbx_altpriority_encoder 2017:10:25:18:06:52:SJ cbx_mgl 2017:10:25:18:08:29:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=8 WIDTHAD=3 data q
--VERSION_BEGIN 17.1 cbx_altpriority_encoder 2017:10:25:18:06:52:SJ cbx_mgl 2017:10:25:18:08:29:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=4 WIDTHAD=2 data q
--VERSION_BEGIN 17.1 cbx_altpriority_encoder 2017:10:25:18:06:52:SJ cbx_mgl 2017:10:25:18:08:29:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=2 WIDTHAD=1 data q
--VERSION_BEGIN 17.1 cbx_altpriority_encoder 2017:10:25:18:06:52:SJ cbx_mgl 2017:10:25:18:08:29:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  ConvIntToFloat_altpriority_encoder_3v7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0)
	 ); 
 END ConvIntToFloat_altpriority_encoder_3v7;

 ARCHITECTURE RTL OF ConvIntToFloat_altpriority_encoder_3v7 IS

 BEGIN

	q(0) <= ( data(1));

 END RTL; --ConvIntToFloat_altpriority_encoder_3v7


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=2 WIDTHAD=1 data q zero
--VERSION_BEGIN 17.1 cbx_altpriority_encoder 2017:10:25:18:06:52:SJ cbx_mgl 2017:10:25:18:08:29:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  ConvIntToFloat_altpriority_encoder_3e8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END ConvIntToFloat_altpriority_encoder_3e8;

 ARCHITECTURE RTL OF ConvIntToFloat_altpriority_encoder_3e8 IS

 BEGIN

	q(0) <= ( data(1));
	zero <= (NOT (data(0) OR data(1)));

 END RTL; --ConvIntToFloat_altpriority_encoder_3e8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  ConvIntToFloat_altpriority_encoder_6v7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0)
	 ); 
 END ConvIntToFloat_altpriority_encoder_6v7;

 ARCHITECTURE RTL OF ConvIntToFloat_altpriority_encoder_6v7 IS

	 SIGNAL  wire_altpriority_encoder10_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_w_lg_w_lg_zero149w150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_w_lg_zero151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_w_lg_zero149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_w_lg_w_lg_zero151w152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_zero	:	STD_LOGIC;
	 COMPONENT  ConvIntToFloat_altpriority_encoder_3v7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  ConvIntToFloat_altpriority_encoder_3e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder11_w_lg_zero149w & wire_altpriority_encoder11_w_lg_w_lg_zero151w152w);
	altpriority_encoder10 :  ConvIntToFloat_altpriority_encoder_3v7
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder10_q
	  );
	wire_altpriority_encoder11_w_lg_w_lg_zero149w150w(0) <= wire_altpriority_encoder11_w_lg_zero149w(0) AND wire_altpriority_encoder11_q(0);
	wire_altpriority_encoder11_w_lg_zero151w(0) <= wire_altpriority_encoder11_zero AND wire_altpriority_encoder10_q(0);
	wire_altpriority_encoder11_w_lg_zero149w(0) <= NOT wire_altpriority_encoder11_zero;
	wire_altpriority_encoder11_w_lg_w_lg_zero151w152w(0) <= wire_altpriority_encoder11_w_lg_zero151w(0) OR wire_altpriority_encoder11_w_lg_w_lg_zero149w150w(0);
	altpriority_encoder11 :  ConvIntToFloat_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder11_q,
		zero => wire_altpriority_encoder11_zero
	  );

 END RTL; --ConvIntToFloat_altpriority_encoder_6v7


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=4 WIDTHAD=2 data q zero
--VERSION_BEGIN 17.1 cbx_altpriority_encoder 2017:10:25:18:06:52:SJ cbx_mgl 2017:10:25:18:08:29:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  ConvIntToFloat_altpriority_encoder_6e8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END ConvIntToFloat_altpriority_encoder_6e8;

 ARCHITECTURE RTL OF ConvIntToFloat_altpriority_encoder_6e8 IS

	 SIGNAL  wire_altpriority_encoder12_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder13_w_lg_w_lg_zero167w168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_w_lg_zero169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_w_lg_zero167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_w_lg_w_lg_zero169w170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_zero	:	STD_LOGIC;
	 COMPONENT  ConvIntToFloat_altpriority_encoder_3e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder13_w_lg_zero167w & wire_altpriority_encoder13_w_lg_w_lg_zero169w170w);
	zero <= (wire_altpriority_encoder12_zero AND wire_altpriority_encoder13_zero);
	altpriority_encoder12 :  ConvIntToFloat_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder12_q,
		zero => wire_altpriority_encoder12_zero
	  );
	wire_altpriority_encoder13_w_lg_w_lg_zero167w168w(0) <= wire_altpriority_encoder13_w_lg_zero167w(0) AND wire_altpriority_encoder13_q(0);
	wire_altpriority_encoder13_w_lg_zero169w(0) <= wire_altpriority_encoder13_zero AND wire_altpriority_encoder12_q(0);
	wire_altpriority_encoder13_w_lg_zero167w(0) <= NOT wire_altpriority_encoder13_zero;
	wire_altpriority_encoder13_w_lg_w_lg_zero169w170w(0) <= wire_altpriority_encoder13_w_lg_zero169w(0) OR wire_altpriority_encoder13_w_lg_w_lg_zero167w168w(0);
	altpriority_encoder13 :  ConvIntToFloat_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder13_q,
		zero => wire_altpriority_encoder13_zero
	  );

 END RTL; --ConvIntToFloat_altpriority_encoder_6e8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  ConvIntToFloat_altpriority_encoder_bv7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0)
	 ); 
 END ConvIntToFloat_altpriority_encoder_bv7;

 ARCHITECTURE RTL OF ConvIntToFloat_altpriority_encoder_bv7 IS

	 SIGNAL  wire_altpriority_encoder8_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder9_w_lg_w_lg_zero140w141w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder9_w_lg_zero142w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder9_w_lg_zero140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder9_w_lg_w_lg_zero142w143w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder9_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder9_zero	:	STD_LOGIC;
	 COMPONENT  ConvIntToFloat_altpriority_encoder_6v7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  ConvIntToFloat_altpriority_encoder_6e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder9_w_lg_zero140w & wire_altpriority_encoder9_w_lg_w_lg_zero142w143w);
	altpriority_encoder8 :  ConvIntToFloat_altpriority_encoder_6v7
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder8_q
	  );
	loop20 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder9_w_lg_w_lg_zero140w141w(i) <= wire_altpriority_encoder9_w_lg_zero140w(0) AND wire_altpriority_encoder9_q(i);
	END GENERATE loop20;
	loop21 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder9_w_lg_zero142w(i) <= wire_altpriority_encoder9_zero AND wire_altpriority_encoder8_q(i);
	END GENERATE loop21;
	wire_altpriority_encoder9_w_lg_zero140w(0) <= NOT wire_altpriority_encoder9_zero;
	loop22 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder9_w_lg_w_lg_zero142w143w(i) <= wire_altpriority_encoder9_w_lg_zero142w(i) OR wire_altpriority_encoder9_w_lg_w_lg_zero140w141w(i);
	END GENERATE loop22;
	altpriority_encoder9 :  ConvIntToFloat_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder9_q,
		zero => wire_altpriority_encoder9_zero
	  );

 END RTL; --ConvIntToFloat_altpriority_encoder_bv7


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=8 WIDTHAD=3 data q zero
--VERSION_BEGIN 17.1 cbx_altpriority_encoder 2017:10:25:18:06:52:SJ cbx_mgl 2017:10:25:18:08:29:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  ConvIntToFloat_altpriority_encoder_be8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END ConvIntToFloat_altpriority_encoder_be8;

 ARCHITECTURE RTL OF ConvIntToFloat_altpriority_encoder_be8 IS

	 SIGNAL  wire_altpriority_encoder14_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder15_w_lg_w_lg_zero177w178w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_w_lg_zero179w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_w_lg_zero177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_w_lg_w_lg_zero179w180w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_zero	:	STD_LOGIC;
	 COMPONENT  ConvIntToFloat_altpriority_encoder_6e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder15_w_lg_zero177w & wire_altpriority_encoder15_w_lg_w_lg_zero179w180w);
	zero <= (wire_altpriority_encoder14_zero AND wire_altpriority_encoder15_zero);
	altpriority_encoder14 :  ConvIntToFloat_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder14_q,
		zero => wire_altpriority_encoder14_zero
	  );
	loop23 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder15_w_lg_w_lg_zero177w178w(i) <= wire_altpriority_encoder15_w_lg_zero177w(0) AND wire_altpriority_encoder15_q(i);
	END GENERATE loop23;
	loop24 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder15_w_lg_zero179w(i) <= wire_altpriority_encoder15_zero AND wire_altpriority_encoder14_q(i);
	END GENERATE loop24;
	wire_altpriority_encoder15_w_lg_zero177w(0) <= NOT wire_altpriority_encoder15_zero;
	loop25 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder15_w_lg_w_lg_zero179w180w(i) <= wire_altpriority_encoder15_w_lg_zero179w(i) OR wire_altpriority_encoder15_w_lg_w_lg_zero177w178w(i);
	END GENERATE loop25;
	altpriority_encoder15 :  ConvIntToFloat_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder15_q,
		zero => wire_altpriority_encoder15_zero
	  );

 END RTL; --ConvIntToFloat_altpriority_encoder_be8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  ConvIntToFloat_altpriority_encoder_rb6 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0)
	 ); 
 END ConvIntToFloat_altpriority_encoder_rb6;

 ARCHITECTURE RTL OF ConvIntToFloat_altpriority_encoder_rb6 IS

	 SIGNAL  wire_altpriority_encoder6_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder7_w_lg_w_lg_zero131w132w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder7_w_lg_zero133w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder7_w_lg_zero131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder7_w_lg_w_lg_zero133w134w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder7_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder7_zero	:	STD_LOGIC;
	 COMPONENT  ConvIntToFloat_altpriority_encoder_bv7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  ConvIntToFloat_altpriority_encoder_be8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder7_w_lg_zero131w & wire_altpriority_encoder7_w_lg_w_lg_zero133w134w);
	altpriority_encoder6 :  ConvIntToFloat_altpriority_encoder_bv7
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder6_q
	  );
	loop26 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder7_w_lg_w_lg_zero131w132w(i) <= wire_altpriority_encoder7_w_lg_zero131w(0) AND wire_altpriority_encoder7_q(i);
	END GENERATE loop26;
	loop27 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder7_w_lg_zero133w(i) <= wire_altpriority_encoder7_zero AND wire_altpriority_encoder6_q(i);
	END GENERATE loop27;
	wire_altpriority_encoder7_w_lg_zero131w(0) <= NOT wire_altpriority_encoder7_zero;
	loop28 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder7_w_lg_w_lg_zero133w134w(i) <= wire_altpriority_encoder7_w_lg_zero133w(i) OR wire_altpriority_encoder7_w_lg_w_lg_zero131w132w(i);
	END GENERATE loop28;
	altpriority_encoder7 :  ConvIntToFloat_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder7_q,
		zero => wire_altpriority_encoder7_zero
	  );

 END RTL; --ConvIntToFloat_altpriority_encoder_rb6

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 2 lpm_compare 1 reg 131 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  ConvIntToFloat_altfp_convert_vpm IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (9 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END ConvIntToFloat_altfp_convert_vpm;

 ARCHITECTURE RTL OF ConvIntToFloat_altfp_convert_vpm IS

	 SIGNAL  wire_altbarrel_shift5_data	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_result	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder2_data	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder2_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL	 exponent_bus_pre_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exponent_bus_pre_reg2	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exponent_bus_pre_reg3	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mag_int_a_reg	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mag_int_a_reg2	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mantissa_pre_round_reg	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 priority_encoder_reg	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 result_reg	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_add_sub1_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_add_sub1_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_add_sub3_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_cmpr4_w_lg_w_lg_alb22w23w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_cmpr4_w_lg_alb21w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_cmpr4_w_lg_alb22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cmpr4_alb	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_max_neg_value_selector18w19w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_sign_int_a5w6w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_max_neg_value_selector17w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_sign_int_a4w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_max_neg_value_selector18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sign_int_a5w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  aclr	:	STD_LOGIC;
	 SIGNAL  bias_value_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  const_bias_value_add_width_int_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exceptions_value :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_bus :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_bus_pre :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_output_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_rounded :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_zero_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  int_a :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  int_a_2s :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  invert_int_a :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  leading_zeroes :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  mag_int_a :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  mantissa_bus :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  mantissa_pre_round :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  mantissa_rounded :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  max_neg_value_selector :	STD_LOGIC;
	 SIGNAL  max_neg_value_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  minus_leading_zero :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  prio_mag_int_a :	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  priority_pad_one_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  shifted_mag_int_a :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  sign_bus :	STD_LOGIC;
	 SIGNAL  sign_int_a :	STD_LOGIC;
	 SIGNAL  zero_padding_w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 COMPONENT  ConvIntToFloat_altbarrel_shift_aof
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clk_en	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(9 DOWNTO 0);
		distance	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		result	:	OUT  STD_LOGIC_VECTOR(9 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  ConvIntToFloat_altpriority_encoder_rb6
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	loop29 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_max_neg_value_selector18w19w(i) <= wire_w_lg_max_neg_value_selector18w(0) AND exponent_zero_w(i);
	END GENERATE loop29;
	loop30 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_sign_int_a5w6w(i) <= wire_w_lg_sign_int_a5w(0) AND int_a(i);
	END GENERATE loop30;
	loop31 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_max_neg_value_selector17w(i) <= max_neg_value_selector AND max_neg_value_w(i);
	END GENERATE loop31;
	loop32 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_sign_int_a4w(i) <= sign_int_a AND int_a_2s(i);
	END GENERATE loop32;
	wire_w_lg_max_neg_value_selector18w(0) <= NOT max_neg_value_selector;
	wire_w_lg_sign_int_a5w(0) <= NOT sign_int_a;
	aclr <= '0';
	bias_value_w <= "01111111";
	clk_en <= '1';
	const_bias_value_add_width_int_w <= "10000111";
	exceptions_value <= (wire_w_lg_w_lg_max_neg_value_selector18w19w OR wire_w_lg_max_neg_value_selector17w);
	exponent_bus <= exponent_rounded;
	exponent_bus_pre <= (wire_cmpr4_w_lg_w_lg_alb22w23w OR wire_cmpr4_w_lg_alb21w);
	exponent_output_w <= wire_add_sub3_result;
	exponent_rounded <= exponent_bus_pre_reg;
	exponent_zero_w <= (OTHERS => '0');
	int_a <= dataa(8 DOWNTO 0);
	int_a_2s <= wire_add_sub1_result;
	invert_int_a <= (NOT int_a);
	leading_zeroes <= (NOT priority_encoder_reg);
	mag_int_a <= (wire_w_lg_w_lg_sign_int_a5w6w OR wire_w_lg_sign_int_a4w);
	mantissa_bus <= mantissa_rounded(22 DOWNTO 0);
	mantissa_pre_round <= ( shifted_mag_int_a(8 DOWNTO 0) & "000000000000000");
	mantissa_rounded <= mantissa_pre_round_reg;
	max_neg_value_selector <= (wire_cmpr4_alb AND sign_int_a_reg2);
	max_neg_value_w <= "10001000";
	minus_leading_zero <= ( zero_padding_w & leading_zeroes);
	prio_mag_int_a <= ( mag_int_a_reg & "1");
	priority_pad_one_w <= (OTHERS => '1');
	result <= result_reg;
	result_w <= ( sign_bus & exponent_bus & mantissa_bus);
	shifted_mag_int_a <= wire_altbarrel_shift5_result(8 DOWNTO 0);
	sign_bus <= sign_int_a_reg5;
	sign_int_a <= dataa(9);
	zero_padding_w <= (OTHERS => '0');
	wire_altbarrel_shift5_data <= ( "0" & mag_int_a_reg2);
	altbarrel_shift5 :  ConvIntToFloat_altbarrel_shift_aof
	  PORT MAP ( 
		aclr => aclr,
		clk_en => clk_en,
		clock => clock,
		data => wire_altbarrel_shift5_data,
		distance => leading_zeroes,
		result => wire_altbarrel_shift5_result
	  );
	wire_altpriority_encoder2_data <= ( prio_mag_int_a & priority_pad_one_w);
	altpriority_encoder2 :  ConvIntToFloat_altpriority_encoder_rb6
	  PORT MAP ( 
		data => wire_altpriority_encoder2_data,
		q => wire_altpriority_encoder2_q
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponent_bus_pre_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponent_bus_pre_reg <= exponent_bus_pre_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponent_bus_pre_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponent_bus_pre_reg2 <= exponent_bus_pre_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponent_bus_pre_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponent_bus_pre_reg3 <= exponent_bus_pre;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mag_int_a_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mag_int_a_reg <= mag_int_a;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mag_int_a_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mag_int_a_reg2 <= mag_int_a_reg;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mantissa_pre_round_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mantissa_pre_round_reg <= mantissa_pre_round;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN priority_encoder_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN priority_encoder_reg <= wire_altpriority_encoder2_q;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN result_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN result_reg <= result_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg1 <= sign_int_a;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg2 <= sign_int_a_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg3 <= sign_int_a_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg4 <= sign_int_a_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg5 <= sign_int_a_reg4;
			END IF;
		END IF;
	END PROCESS;
	wire_add_sub1_datab <= "000000001";
	add_sub1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 9,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => invert_int_a,
		datab => wire_add_sub1_datab,
		result => wire_add_sub1_result
	  );
	add_sub3 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_WIDTH => 8,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => const_bias_value_add_width_int_w,
		datab => minus_leading_zero,
		result => wire_add_sub3_result
	  );
	loop33 : FOR i IN 0 TO 7 GENERATE 
		wire_cmpr4_w_lg_w_lg_alb22w23w(i) <= wire_cmpr4_w_lg_alb22w(0) AND exponent_output_w(i);
	END GENERATE loop33;
	loop34 : FOR i IN 0 TO 7 GENERATE 
		wire_cmpr4_w_lg_alb21w(i) <= wire_cmpr4_alb AND exceptions_value(i);
	END GENERATE loop34;
	wire_cmpr4_w_lg_alb22w(0) <= NOT wire_cmpr4_alb;
	cmpr4 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		alb => wire_cmpr4_alb,
		dataa => exponent_output_w,
		datab => bias_value_w
	  );

 END RTL; --ConvIntToFloat_altfp_convert_vpm
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ConvIntToFloat IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		dataa		: IN STD_LOGIC_VECTOR (9 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END ConvIntToFloat;


ARCHITECTURE RTL OF convinttofloat IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (31 DOWNTO 0);



	COMPONENT ConvIntToFloat_altfp_convert_vpm
	PORT (
			clock	: IN STD_LOGIC ;
			dataa	: IN STD_LOGIC_VECTOR (9 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(31 DOWNTO 0);

	ConvIntToFloat_altfp_convert_vpm_component : ConvIntToFloat_altfp_convert_vpm
	PORT MAP (
		clock => clock,
		dataa => dataa,
		result => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altfp_convert"
-- Retrieval info: CONSTANT: OPERATION STRING "INT2FLOAT"
-- Retrieval info: CONSTANT: ROUNDING STRING "TO_NEAREST"
-- Retrieval info: CONSTANT: WIDTH_DATA NUMERIC "10"
-- Retrieval info: CONSTANT: WIDTH_EXP_INPUT NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_EXP_OUTPUT NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_INT NUMERIC "10"
-- Retrieval info: CONSTANT: WIDTH_MAN_INPUT NUMERIC "23"
-- Retrieval info: CONSTANT: WIDTH_MAN_OUTPUT NUMERIC "23"
-- Retrieval info: CONSTANT: WIDTH_RESULT NUMERIC "32"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: USED_PORT: dataa 0 0 10 0 INPUT NODEFVAL "dataa[9..0]"
-- Retrieval info: CONNECT: @dataa 0 0 10 0 dataa 0 0 10 0
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL ConvIntToFloat.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ConvIntToFloat.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ConvIntToFloat.bsf TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ConvIntToFloat_inst.vhd TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ConvIntToFloat.inc TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ConvIntToFloat.cmp TRUE TRUE
-- Retrieval info: LIB_FILE: lpm
