CompPWM_inst : CompPWM PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		alb	 => alb_sig
	);
