ConstSigma_inst : ConstSigma PORT MAP (
		result	 => result_sig
	);
