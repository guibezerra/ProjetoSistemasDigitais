Comparador_somador_inst : Comparador_somador PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		aneb	 => aneb_sig
	);
