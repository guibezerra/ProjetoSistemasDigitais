Contator_Somador_inst : Contator_Somador PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
