Constantes_inst : Constantes PORT MAP (
		result	 => result_sig
	);
