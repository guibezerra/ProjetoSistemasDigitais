ContadorPWM_inst : ContadorPWM PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
