constante_255_inst : constante_255 PORT MAP (
		result	 => result_sig
	);
